`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/08/2022 02:40:33 PM
// Design Name: 
// Module Name: imgen
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module imgen;
reg [31:0] inst_out;
wire  [31:0] immgenout;
reg clk,rst;

immgen ig1 (.instr(inst_out),.out(immgenout),.clk(clk),.rst(rst));

initial
begin
clk=0;
rst=0;
inst_out=32'b01111010101011000110001000000011;
#10;
clk=1;
rst=0;
inst_out=32'b01111010101011000110001000000011;
#10;
clk=0;
rst=1;
inst_out=32'b01111010101011000110001000000011;
#10;
clk=1;
rst=1;
inst_out=32'b01111010101011000110001000000011;
#10;
/////
clk=0;
rst=0;
inst_out=32'b10111010111010011000101000100011;
#10;
clk=1;
rst=0;
inst_out=32'b10111010111010011000101000100011 ;
#10;
clk=0;
rst=1;
inst_out=32'b10111010111010011000101000100011 ;
#10;
clk=1;
rst=1;
inst_out=32'b10111010111010011000101000100011 ;
#10;
////////////////
clk=0;
rst=0;
inst_out=32'b01100111000110011110000001100011;
#10;
clk=1;
rst=0;
inst_out=32'b01100111000110011110000001100011 ;
#10;
clk=0;
rst=1;
inst_out=32'b01100111000110011110000001100011 ;
#10;
clk=1;
rst=1;
inst_out=32'b01100111000110011110000001100011 ;
#10;
////////////
clk=0;
rst=0;
inst_out=32'b11111111000111100001100000010011;
#10;
clk=1;
rst=0;
inst_out=32'b11111111000111100001100000010011 ;
#10;
clk=0;
rst=1;
inst_out=32'b11111111000111100001100000010011 ;
#10;
clk=1;
rst=1;
inst_out=32'b11111111000111100001100000010011 ;
#10;
////////////
clk=0;
rst=0;
inst_out=32'b11111111110000001100000001100111;
#10;
clk=1;
rst=0;
inst_out=32'b11111111110000001100000001100111 ;
#10;
clk=0;
rst=1;
inst_out=32'b11111111110000001100000001100111 ;
#10;
clk=1;
rst=1;
inst_out=32'b11111111110000001100000001100111 ;
#10;
////////
clk=0;
rst=0;
inst_out=32'b00001111111111111100000001101111;
#10;
clk=1;
rst=0;
inst_out=32'b00001111111111111100000001101111 ;
#10;
clk=0;
rst=1;
inst_out=32'b00001111111111111100000001101111 ;
#10;
clk=1;
rst=1;
inst_out=32'b00001111111111111100000001101111 ;
end


endmodule
